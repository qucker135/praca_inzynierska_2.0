----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 21.12.2022 11:52:24
-- Design Name: 
-- Module Name: program_memory - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity program_memory is
    Port ( clk : in STD_LOGIC;
           addr_in : in STD_LOGIC_VECTOR (10 downto 0);
           dout : out STD_LOGIC_VECTOR (13 downto 0));
end program_memory;

architecture Behavioral of program_memory is

    type program_memory_type is array (0 to 2047) of STD_LOGIC_VECTOR(13 downto 0);
    
    signal mem_contents : program_memory_type := (
        0 => B"00_1111_1111_1111", -- INCFSZ
        1 => B"00_1111_1111_1111", -- INCFSZ
        2 => B"00_1111_1111_1111", -- INCFSZ
        3 => B"00_1011_1111_1111", -- DECFSZ
        4 => B"00_1011_1111_1111", -- DECFSZ
        5 => B"00_1011_1111_1111", -- DECFSZ
        6 => B"00_1011_1111_1111", -- DECFSZ
        7 => B"00_1011_1111_1111", -- DECFSZ
        8 => B"00_1111_1111_1111", -- INCFSZ
        9 => B"00_1111_1111_1111", -- INCFSZ
       10 => B"00_1111_1111_1111", -- INCFSZ
       11 => B"00_1111_1111_1111", -- INCFSZ
       12 => B"00_1111_1111_1111", -- INCFSZ
       13 => B"00_1011_1111_1111", -- DECFSZ
       14 => B"00_1011_1111_1111", -- DECFSZ
       15 => B"00_1011_1111_1111", -- DECFSZ
       16 => B"00_1011_1111_1111", -- DECFSZ
       17 => B"00_1011_1111_1111", -- DECFSZ
       18 => B"00_1111_1111_1111", -- INCFSZ
       19 => B"00_1111_1111_1111", -- INCFSZ
       20 => B"00_1111_1111_1111", -- INCFSZ
       21 => B"00_1111_1111_1111", -- INCFSZ
       22 => B"00_1111_1111_1111", -- INCFSZ
        others => B"00_0000_0000_0000");

begin

    process(clk)
    begin
        if rising_edge(clk) then
            dout <= mem_contents(to_integer(unsigned(addr_in)));
        end if;
    end process;

end Behavioral;
